
package pkg1;
    function int f1(int x);
        return `ADD(x, 5);
    endfunction
endpackage

`define UNUSED_WIRE(name) wire name; assign name = 1'b0;

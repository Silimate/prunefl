module mylib1;
endmodule


module c();
  d d_mod();
endmodule

module a();
  b b_mod();
endmodule

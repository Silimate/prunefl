
  module top_module(input [a_pkg::a_param - 1:0] in, output [a_pkg::a_param - 1:0] out);
    assign out = ~in;
  endmodule
  

`define MODULE_B_NAME module_b

module utils #(parameter DEPTH = 4) (
    input wire in,
    output wire out
);
    assign out = in;
endmodule


  package b_pkg;
    localparam int b_param = 1;
  endpackage
  


  package a_pkg;
    localparam int a_param = b_pkg::b_param;
  endpackage
  

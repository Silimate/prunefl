`include "macros.vh"

module `MODULE_B_NAME (
    input wire clk,
    input wire in_b,
    output wire out_b
);
    assign out_b = in_b;
endmodule

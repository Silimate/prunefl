
`define ADD(x, y) ((x) + (y))
`define MUL(x, y) ((x) * (y))
`define MACRO_FUNC `ADD(`MUL(2, 3), 4)

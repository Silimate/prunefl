function void Misc::sayHi(string target);
  $display("Hi, %s!", target);
endfunction

module dummy();

endmodule

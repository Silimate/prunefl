`define DEFAULT_WIDTH 8
`define CONNECT(a, b) assign a = b
`include "macros.vh" // TODO: Handle explicit include
`define LITERALLY_USELESS `UNUSED_WIRE(useless)
`define CORE_LOGIC_NAME core_logic

module top_module;
  alu u_alu();
  mylib1 u1();
endmodule

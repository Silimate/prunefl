

module d();
  initial $display("hi");
endmodule

module b();
  c c_cmod();
endmodule

module top_module();
  a a_mod();
endmodule

module mylib2;
endmodule

class Misc;
  extern function void sayHi(string target);
endclass
